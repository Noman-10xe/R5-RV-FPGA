B8201073B0201073
0000011300000093
0000021300000193
0000031300000293
0000041300000393
0000051300000493
0000061300000593
0000071300000693
0000081300000793
0000091300000893
00000A1300000993
00000B1300000A93
00000C1300000B93
00000D1300000C93
00000E1300000D93
00000F1300000E93
5555533700000F93
7C03107355530313
0701819300003197
8681011300004117
8605051300003517
8585859300003597
0005202300B57863
FEB56CE300450513
00000513634000EF
00C000EF00000593
000000000000006F
00100793FC010113
0001041302812C23
02112E2300F12223
0321282302912A23
0281069300012023
0007A70300040793
004787930047A603
00E7A22300C70733
248000EFFED796E3
8A45051300001537
03040493570000EF
0004258300001937
004404138C490513
FE8498E3558000EF
000507930000006F
000716630007C703
0000806740A78533
FEDFF06F00178793
00812423FF010113
00A0079300112623
00F5166300050413
FE5FF0EF00D00513
0147278380002737
FE078CE30207F793
00C1208300872023
0000051300812403
0000806701010113
040786630105A783
FF01011304050463
0005A48300912223
0011262300812423
0044278300058413
00C4450300F4DA63
F85FF0EF00148493
00C12083FEDFF06F
0041248300812403
0000806701010113
F901011300008067
0005899305312E23
06812423000015B7
8C85859306912223
0006049300050413
0110061300810513
0721202306112623
000015B7550000EF
8DC5859301100613
53C000EF01C10513
0CF9946300A00793
408005330C045263
0184A78300100613
0007946300810713
0301091301C10713
0009079300A00693
0AD9986300F00593
0090081300A00593
0017879302B576B3
0006C68300D706B3
02B556B3FED78FA3
0006086308A86063
00E7802302D00713
0007802300178793
FFF7841300090513
00A4A023E85FF0EF
000485930144A503
0015351300040993
01246863ED1FF0EF
408987B301C4A703
0144A50306E7C263
EB5FF0EF00048593
0681240306C12083
0601290306412483
0701011305C12983
0004051300008067
F41FF06F00000613
F65FF06F00068513
00F5769300068513
0006C68300D706B3
FED78FA300178793
FEA5E2E300455693
FFF40413F5DFF06F
E0DFF0EF00144503
800027B7F85FF06F
00E7AA230FF00713
00E7A62308000713
00E7A02301B00713
00E7A62300300713
00E7A42308700713
000080670007A223
F901011300008737
06812423FFF70793
05512A2305412C23
0611262305A12023
0721202306912223
0561282305312E23
0581242305712623
03B12E2305912223
00058D1300050413
00F1262302500A13
0004450306400A93
06C1208304051063
0641248306812403
05C1298306012903
05412A8305812A03
04C12B8305012B03
04412C8304812C03
03C12D8304012D03
0000806707010113
D35FF0EF01450663
00C127831140006F
00E10E2302000713
0201202300A00713
00F12C2302012223
0004049302E12623
0090099300000B13
00100C1307300B93
05C00D9302E00C93
001404130014C503
0FF77713FD050713
040B026308E9E463
00A0059300000713
00100B1301C0006F
FD5FF06F00040493
0014041302B70733
0004468300E68733
0FF6F613FD068693
00E12C23FEC9F4E3
FD5FF06FFFF40413
00E5146303000713
0000071300A10E23
0004468300A00593
0FF6F613FD068693
00E12A2300C9F863
FCDFF06F03812023
0014041302B70733
FD9FF06F00E68733
0FF6F693FBF50693
02C1242301A6B613
0005071301900793
0205071300D7E463
02EACE6309570863
00ECCC63F79702E3
02D0069307470863
0014041306D70863
0FB70A63E9DFF06F
FED718E306300693
004D0493000D4503
0680006FC01FF0EF
02EBC66307770663
F2F702E306C00793
FCD714E307000693
004D049300800713
0101061302E12623
0300006F01000593
00D70E6307500693
FD9FF06F07800693
E81FF06F02500513
EE5FF06F03812223
01010613004D0493
000D250300A00593
00048D13C35FF0EF
000D2483F75FF06F
00048513004D0913
00A12823B65FF0EF
0101059302412503
BB5FF0EF00153513
020792630004C783
B41FF0EF00048513
0241250300A12823
00090D1301010593
F29FF06FB91FF0EF
FFF7871301812783
FC078AE300E12C23
FFF4C50300148493
FBDFF06FB29FF0EF
02E50E6306800713
0610071300A76C63
B0DFF0EF02E50463
E3DFF06F00248413
02E5026306E00713
FEE514E307200713
FE1FF06F00D00513
FD9FF06F00700513
FD1FF06F00800513
FC9FF06F00A00513
00812C23FC010113
02B1222300112E23
02D1262302C12423
02F12A2302E12823
03112E2303012C23
00050A6300000413
00B1262302410593
00050413CC9FF0EF
A8DFF0EF00A00513
01C1208300040513
0401011301812403
FF01011300008067
0121202300812423
9004041300000417
8F89091300000917
0011262340890933
4029591300912223
0000049300090E63
0014849300042783
000780E700440413
00000417FE9918E3
000009178C440413
408909338BC90913
00090E6340295913
0004278300000493
0044041300148493
FE9918E3000780E7
0081240300C12083
0001290300412483
0000806701010113
0037F79300A5C7B3
0607926300C508B3
04C7FE6300300793
0005071300357793
FFC8F61306079863
08F76C63FE060793
0005869302C77C63
0006A80300070793
0046869300478793
FEC7E8E3FF07AE23
40E787B3FFF60793
00478793FFC7F793
00F585B300F70733
0000806701176863
FF157CE300050713
001707130005C783
FEF70FA300158593
00008067FF1768E3
001707130005C683
FED70FA300377793
F80780E300158593
001707130005C683
FED70FA300377793
FC079AE300158593
0005A683F65FF06F
0085AF830045A283
0105AE8300C5AF03
0185A3030145AE03
0245859301C5A803
FFC5A68300D72023
01F7242300572223
01D7282301E72623
00672C2301C72A23
0247071301072E23
FAF768E3FED72E23
6F626946F19FF06F
655320696363616E
6946282073656972
3A29323120747372
000064250000000A
3736353433323130
4645444342413938
3332313000000000
6261393837363534
0000000066656463
0000000000000000
