B8201073B0201073
0000011300000093
0000021300000193
0000031300000293
0000041300000393
0000051300000493
0000061300000593
0000071300000693
0000081300000793
0000091300000893
00000A1300000993
00000B1300000A93
00000C1300000B93
00000D1300000C93
00000E1300000D93
00000F1300000E93
5555533700000F93
7C03107355530313
9181819300003197
1101011300003117
1085051300002517
1005859300002597
0005202300B57863
FEB56CE300450513
00000513048000EF
00C000EF00000593
000000000000006F
80001737000107B7
40F72423FFF78793
4006A703800016B7
00F7F79301075793
00E787B301C75713
FE9FF06F40F6A223
00812423FF010113
0000041701212023
00000917EEC40413
40890933EE490913
0091222300112623
00090E6340295913
0004278300000493
0044041300148493
FE9918E3000780E7
EB04041300000417
EA89091300000917
4029591340890933
0000049300090E63
0014849300042783
000780E700440413
00C12083FE9918E3
0041248300812403
0101011300012903
0000000000008067
