B8201073B0201073
0000011300000093
0000021300000193
0000031300000293
0000041300000393
0000051300000493
0000061300000593
0000071300000693
0000081300000793
0000091300000893
00000A1300000993
00000B1300000A93
00000C1300000B93
00000D1300000C93
00000E1300000D93
00000F1300000E93
5555533700000F93
7C03107355530313
9701819300003197
1681011300003117
1605051300002517
1585859300002597
0005202300B57863
FEB56CE300450513
0000051309C000EF
00C000EF00000593
000000000000006F
00812423FF010113
8000173700112623
02F72C230F000793
FFF78793000107B7
8000143740F72423
0C80051340042783
02F42E234107D793
FEDFF06F008000EF
00012423FF010113
00A7C66300812783
0000806701010113
00C1278300012623
0081278300F05A63
00F1242300178793
00C12783FD9FF06F
00F1262300178793
FF010113FDDFF06F
0121202300812423
E984041300000417
E909091300000917
0011262340890933
4029591300912223
0000049300090E63
0014849300042783
000780E700440413
00000417FE9918E3
00000917E5C40413
40890933E5490913
00090E6340295913
0004278300000493
0044041300148493
FE9918E3000780E7
0081240300C12083
0001290300412483
0000806701010113
0000000000000000
