B8201073B0201073
0000011300000093
0000021300000193
0000031300000293
0000041300000393
0000051300000493
0000061300000593
0000071300000693
0000081300000793
0000091300000893
00000A1300000993
00000B1300000A93
00000C1300000B93
00000D1300000C93
00000E1300000D93
00000F1300000E93
5555533700000F93
7C03107355530313
9901819300003197
1881011300003117
1805051300002517
1785859300002597
0005202300B57863
FEB56CE300450513
000005130BC000EF
050000EF00000593
000000000000006F
00112023FF810113
0005041300812223
0010039300000293
000003130082DE63
0013031300735663
00128293FF9FF06F
00012083FE9FF06F
0081011300412403
FF41011300008067
0081222300112023
8000143700912423
800014B740040413
000102B703848493
00542423FFF28293
0054A0230F000293
0102D29300042283
0C8005130054A223
FEDFF06FF79FF0EF
0041240300012083
00C1011300812483
FF01011300008067
0121202300812423
E784041300000417
E709091300000917
0011262340890933
4029591300912223
0000049300090E63
0014849300042783
000780E700440413
00000417FE9918E3
00000917E3C40413
40890933E3490913
00090E6340295913
0004278300000493
0044041300148493
FE9918E3000780E7
0081240300C12083
0001290300412483
0000806701010113
0000000000000000
