B8201073B0201073
0000011300000093
0000021300000193
0000031300000293
0000041300000393
0000051300000493
0000061300000593
0000071300000693
0000081300000793
0000091300000893
00000A1300000993
00000B1300000A93
00000C1300000B93
00000D1300000C93
00000E1300000D93
00000F1300000E93
5555533700000F93
7C03107355530313
0B81819300003197
8B01011300004117
8A85051300003517
8A05859300003597
0005202300B57863
FEB56CE300450513
00000513660000EF
00C000EF00000593
000000000000006F
000015B7FC010113
8D05859303000613
02112E2300010513
02912A2302812C23
6B8000EF03212823
038000EF00010513
00001537288000EF
5B0000EF90050513
0301049300010413
0004258300001937
0044041391090513
FE9418E3594000EF
00B007130000006F
0000069300050793
0007A6030200006F
00C5D6630047A583
00C7A22300B7A023
0047879300168693
FFF70713FEE6C2E3
00008067FC0718E3
0007C70300050793
40A7853300071663
0017879300008067
FF010113FEDFF06F
0011262300812423
0005041300A00793
00D0051300F51663
80002737FE5FF0EF
0207F79301472783
00872023FE078CE3
0081240300C12083
0101011300000513
0105A78300008067
0405046304078663
00912223FF010113
008124230005A483
0005841300112623
00F4DA6300442783
0014849300C44503
FEDFF06FF85FF0EF
0081240300C12083
0101011300412483
0000806700008067
05312E23F9010113
000015B700058993
0691222306812423
0005041391458593
0081051300060493
0611262301100613
550000EF07212023
01100613000015B7
01C1051392858593
00A0079353C000EF
0C0452630CF99463
0010061340800533
008107130184A783
01C1071300079463
00A0069303010913
00F0059300090793
00A005930AD99863
02B576B300900813
00D706B300178793
FED78FA30006C683
08A8606302B556B3
02D0071300060863
0017879300E78023
0009051300078023
E85FF0EFFFF78413
0144A50300A4A023
0004099300048593
ED1FF0EF00153513
01C4A70301246863
06E7C263408987B3
000485930144A503
06C12083EB5FF0EF
0641248306812403
05C1298306012903
0000806707010113
0000061300040513
00068513F41FF06F
00068513F65FF06F
00D706B300F57693
001787930006C683
00455693FED78FA3
F5DFF06FFEA5E2E3
00144503FFF40413
F85FF06FE0DFF0EF
0FF00713800027B7
0800071300E7AA23
01B0071300E7A623
0030071300E7A023
0870071300E7A623
0007A22300E7A423
0000873700008067
FFF70793F9010113
05412C2306812423
05A1202305512A23
0691222306112623
05312E2307212023
0571262305612823
0591222305812423
0005041303B12E23
02500A1300058D13
06400A9300F12623
0405106300044503
0681240306C12083
0601290306412483
05812A0305C12983
05012B0305412A83
04812C0304C12B83
04012D0304412C83
0701011303C12D83
0145066300008067
1140006FD35FF0EF
0200071300C12783
00A0071300E10E23
0201222302012023
02E1262300F12C23
00000B1300040493
07300B9300900993
02E00C9300100C13
0014C50305C00D93
FD05071300140413
08E9E4630FF77713
00000713040B0263
01C0006F00A00593
0004049300100B13
02B70733FD5FF06F
00E6873300140413
FD06869300044683
FEC9F4E30FF6F613
FFF4041300E12C23
03000713FD5FF06F
00A10E2300E51463
00A0059300000713
FD06869300044683
00C9F8630FF6F613
0381202300E12A23
02B70733FCDFF06F
00E6873300140413
FBF50693FD9FF06F
01A6B6130FF6F693
0190079302C12423
00D7E46300050713
0957086302050713
F79702E302EACE63
0747086300ECCC63
06D7086302D00693
E9DFF06F00140413
063006930FB70A63
000D4503FED718E3
C01FF0EF004D0493
077706630680006F
06C0079302EBC663
07000693F2F702E3
00800713FCD714E3
02E12623004D0493
0100059301010613
075006930300006F
0780069300D70E63
02500513FD9FF06F
03812223E81FF06F
004D0493EE5FF06F
00A0059301010613
C35FF0EF000D2503
F75FF06F00048D13
004D0913000D2483
B65FF0EF00048513
0241250300A12823
0015351301010593
0004C783BB5FF0EF
0004851302079263
00A12823B41FF0EF
0101059302412503
B91FF0EF00090D13
01812783F29FF06F
00E12C23FFF78713
00148493FC078AE3
B29FF0EFFFF4C503
06800713FBDFF06F
00A76C6302E50E63
02E5046306100713
00248413B0DFF0EF
06E00713E3DFF06F
0720071302E50263
00D00513FEE514E3
00700513FE1FF06F
00800513FD9FF06F
00A00513FD1FF06F
FC010113FC9FF06F
00112E2300812C23
02C1242302B12223
02E1282302D12623
03012C2302F12A23
0000041303112E23
0241059300050A63
CC9FF0EF00B12623
00A0051300050413
00040513A8DFF0EF
0181240301C12083
0000806704010113
00812423FF010113
0000041701212023
000009178D440413
408909338CC90913
0091222300112623
00090E6340295913
0004278300000493
0044041300148493
FE9918E3000780E7
8984041300000417
8909091300000917
4029591340890933
0000049300090E63
0014849300042783
000780E700440413
00C12083FE9918E3
0041248300812403
0101011300012903
00A5C7B300008067
00C508B30037F793
0030079306079263
0035779304C7FE63
0607986300050713
FE060793FFC8F613
02C77C6308F76C63
0007079300058693
004787930006A803
FF07AE2300468693
FFF60793FEC7E8E3
FFC7F79340E787B3
00F7073300478793
0117686300F585B3
0005071300008067
0005C783FF157CE3
0015859300170713
FF1768E3FEF70FA3
0005C68300008067
0037779300170713
00158593FED70FA3
0005C683F80780E3
0037779300170713
00158593FED70FA3
F65FF06FFC079AE3
0045A2830005A683
00C5AF030085AF83
0145AE030105AE83
01C5A8030185A303
00D7202302458593
00572223FFC5A683
01E7262301F72423
01C72A2301D72823
01072E2300672C23
FED72E2302470713
F19FF06FFAF768E3
FFFFFFFE0000000D
000003D600000003
0000007900000021
00000049000001E2
000000650000005E
0000000A00000013
6120646574726F53
0000003A79617272
3332313000006425
4241393837363534
0000000046454443
3736353433323130
6665646362613938
0000000000000000
